library ieee;
use ieee.std_logic_1164.all;

package CHAR_LIB is
    constant A      : std_logic_vector(7 downto 0) := x"41";
    constant B      : std_logic_vector(7 downto 0) := x"42";
    constant C      : std_logic_vector(7 downto 0) := x"43";
    constant D      : std_logic_vector(7 downto 0) := x"44";
    constant E      : std_logic_vector(7 downto 0) := x"45";
    constant F      : std_logic_vector(7 downto 0) := x"46";
    constant G      : std_logic_vector(7 downto 0) := x"47";
    constant H      : std_logic_vector(7 downto 0) := x"48";
    constant I      : std_logic_vector(7 downto 0) := x"49";
    constant J      : std_logic_vector(7 downto 0) := x"4A";
    constant K      : std_logic_vector(7 downto 0) := x"4B";
    constant L      : std_logic_vector(7 downto 0) := x"4C";
    constant M      : std_logic_vector(7 downto 0) := x"4D";
    constant N      : std_logic_vector(7 downto 0) := x"4E";
    constant O      : std_logic_vector(7 downto 0) := x"4F";
    constant P      : std_logic_vector(7 downto 0) := x"50";
    constant Q      : std_logic_vector(7 downto 0) := x"51";
    constant R      : std_logic_vector(7 downto 0) := x"52";
    constant S      : std_logic_vector(7 downto 0) := x"53";
    constant T      : std_logic_vector(7 downto 0) := x"54";
    constant U      : std_logic_vector(7 downto 0) := x"55";
    constant V      : std_logic_vector(7 downto 0) := x"56";
    constant W      : std_logic_vector(7 downto 0) := x"57";
    constant X      : std_logic_vector(7 downto 0) := x"58";
    constant Y      : std_logic_vector(7 downto 0) := x"59";
    constant Z      : std_logic_vector(7 downto 0) := x"5A";

    constant SPACE  : std_logic_vector(7 downto 0) := x"20";
    constant COLON  : std_logic_vector(7 downto 0) := x"3A";
    constant ARROW  : std_logic_vector(7 downto 0) := x"1B";
    constant LESS_THAN  : std_logic_vector(7 downto 0) := x"3c";
    constant DASH   : std_logic_vector(7 downto 0) := x"2D";

    constant a_l    : std_logic_vector(7 downto 0) := x"61";
    constant b_l    : std_logic_vector(7 downto 0) := x"62";
    constant c_l    : std_logic_vector(7 downto 0) := x"63";
    constant d_l    : std_logic_vector(7 downto 0) := x"64";
    constant e_l    : std_logic_vector(7 downto 0) := x"65";
    constant f_l    : std_logic_vector(7 downto 0) := x"66";
    constant g_l    : std_logic_vector(7 downto 0) := x"67";
    constant h_l    : std_logic_vector(7 downto 0) := x"68";
    constant i_l    : std_logic_vector(7 downto 0) := x"69";
    constant j_l    : std_logic_vector(7 downto 0) := x"6A";
    constant k_l    : std_logic_vector(7 downto 0) := x"6B";
    constant l_l    : std_logic_vector(7 downto 0) := x"6C";
    constant m_l    : std_logic_vector(7 downto 0) := x"6D";
    constant n_l    : std_logic_vector(7 downto 0) := x"6E";
    constant o_l    : std_logic_vector(7 downto 0) := x"6F";
    constant p_l    : std_logic_vector(7 downto 0) := x"70";
    constant q_l    : std_logic_vector(7 downto 0) := x"71";
    constant r_l    : std_logic_vector(7 downto 0) := x"72";
    constant s_l    : std_logic_vector(7 downto 0) := x"73";
    constant t_l    : std_logic_vector(7 downto 0) := x"74";
    constant u_l    : std_logic_vector(7 downto 0) := x"75";
    constant v_l    : std_logic_vector(7 downto 0) := x"76";
    constant w_l    : std_logic_vector(7 downto 0) := x"77";
    constant x_l    : std_logic_vector(7 downto 0) := x"78";
    constant y_l    : std_logic_vector(7 downto 0) := x"79";
    constant z_l    : std_logic_vector(7 downto 0) := x"7A";

    constant char_0 : std_logic_vector(7 downto 0) := x"30";
    constant char_1 : std_logic_vector(7 downto 0) := x"31";
    constant char_2 : std_logic_vector(7 downto 0) := x"32";
    constant char_3 : std_logic_vector(7 downto 0) := x"33";
    constant char_4 : std_logic_vector(7 downto 0) := x"34";
    constant char_5 : std_logic_vector(7 downto 0) := x"35";
    constant char_6 : std_logic_vector(7 downto 0) := x"36";
    constant char_7 : std_logic_vector(7 downto 0) := x"37";
    constant char_8 : std_logic_vector(7 downto 0) := x"38";
    constant char_9 : std_logic_vector(7 downto 0) := x"39";

end CHAR_LIB;
