doodle_boy_logo_inst : doodle_boy_logo PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
